** Profile: "SCHEMATIC1-test"  [ C:\Repos\LSG-Microcontroller-EMobility\CellBatteryHealthyCheck\orcad tests\zener_best_practices-pspicefiles\schematic1\test.sim ] 

** Creating circuit file "test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../zener_best_practices-pspicefiles/zener_best_practices.lib" 
* From [PSPICE NETLIST] section of C:\Users\luigi.santagada\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 5 0 0.001 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
